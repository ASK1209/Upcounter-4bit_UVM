package up_counter_pkg;
	import uvm_pkg::*;
	`include "uvm_macros.svh"
	`include "up_xtn.sv"
	`include "up_config.sv"
	`include "up_sequencer.sv"
	`include "up_driver.sv"
	`include "up_monitor.sv"
	`include "up_seqs.sv"
	`include "up_agent.sv"
	`include "up_ref_model.sv"
	`include "up_scoreboard.sv"
	`include "up_env.sv"
	`include "up_test.sv"
endpackage
